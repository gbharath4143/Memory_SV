class bfm_mem();
	task run();		
		$display("BFM");
	endtask
endclass
