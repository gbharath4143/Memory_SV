class coverage_mem();
	task run();		
		$display("COV");
	endtask
endclass
