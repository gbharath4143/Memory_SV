class scoreboard_mem();
	task run();		
		$display("SBD");
	endtask
endclass
