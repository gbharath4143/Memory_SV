class monitor_mem();
	task run();		
		$display("Monitor");
	endtask
endclass
