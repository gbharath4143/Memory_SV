`include "common_mem.sv"
`include "interface_mem.sv"
`include "txn_mem.sv"

`include "coverage_mem.sv"
`include "scoreboard_mem.sv"
`include "monitor_mem.sv"
`include "bfm_mem.sv"
`include "generator_mem.sv"

`include "agent_mem.sv"
`include "env_mem.sv"
`include "top_mem.sv"

`include "memory.sv"
